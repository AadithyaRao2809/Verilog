`include "alu.v"
`include "register.v"

module reg_alu()